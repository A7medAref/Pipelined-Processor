module moduleName ();
    
endmodule